module xor2_tb(); 

