module an2_tb(); 

an2 andtemp();
initial
begin
end
endmodule
