module and2_tb(); 

 reg a,b;

 wire  c;

and2 andtemp();
initial
begin
end
endmodule
